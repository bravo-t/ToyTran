Vin 3 0 pwl(
  0 0 
  1ns 5)
R2 3 2 1000
R1 1 0 1000
C1 1 0 1E-6
C2 2 1 10E-6
L1 1 0 0.001

.tran 1ps 10ns