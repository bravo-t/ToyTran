VVDD Pos Gnd 5V
LInd1 Pos IndOut 1
CCap1 IndOut Gnd 1u

.tran 100us 100ms
.option method=gear2
.plot tran V(IndOut)
.debug 0
