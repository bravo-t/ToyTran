Vg 1 0 4
Vx 3 2 6
R1 1 2 1
R2 2 0 4
R3 3 0 2
It 1 2 1

.tran 1ns 100ns