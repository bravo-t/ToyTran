VVDD POS GND 5
RRes1 POS ResOUT 1k
CCap2 ResOUT GND 1u
*RRes2 3 4 1k
*RRes3 4 0 1k

.tran 1us 10us
*.option method=gear2
.option method=trap
*.plot tran V(2) V(0) V(1) I(Res1) I(Cap2) I(VDD)
.plot tran V(ResOUT) 
.debug 1
