V1 1 0 12
R1 1 2 1000
R2 2 0 2000
R3 2 0 2000

.tran 1ns 1000ns
.debug 0